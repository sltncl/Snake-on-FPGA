LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

-- Define the snake_pkg package
PACKAGE snake_pkg IS

	-- Display and game area dimensions
	CONSTANT display_width  : INTEGER := 1368;  -- Display width in pixels
   CONSTANT display_height : INTEGER := 768;   -- Display height in pixels
   CONSTANT game_width     : INTEGER := 930;   -- Game area width in pixels
   CONSTANT game_height    : INTEGER := 620;   -- Game area height in pixels
	
	-- Snake configuration
   CONSTANT max_snake_length 	: INTEGER := 32;  -- Maximum number of snake segments
   CONSTANT rect_width  		: INTEGER := 31;       -- Width of each snake segment block
   CONSTANT rect_height 		: INTEGER := 31;       -- Height of each snake segment block
	
	-- Game area boundary coordinates
   CONSTANT game_left   : INTEGER := (display_width - game_width) / 2; -- Left coordinate of the game area
   CONSTANT game_right  : INTEGER := game_left + game_width;           -- Right coordinate of the game area
   CONSTANT game_top    : INTEGER := (display_height - game_height) / 2; -- Top coordinate of the game area
   CONSTANT game_bottom : INTEGER := game_top + game_height;           -- Bottom coordinate of the game area

	-- Type declarations for the snake and images
	TYPE snake_segment IS RECORD
		x : INTEGER;
      y : INTEGER;
   END RECORD;	
	
	TYPE snake_array IS ARRAY (0 TO max_snake_length - 1) OF snake_segment;
	TYPE image_type IS ARRAY (0 TO 30, 0 TO 30) OF STD_LOGIC_VECTOR(11 DOWNTO 0);
	TYPE score_image_type IS ARRAY (0 TO 30, 0 TO 185) OF STD_LOGIC_VECTOR(11 DOWNTO 0); 
	TYPE gameOver_image_type IS ARRAY (0 TO 39, 0 TO 367) OF STD_LOGIC_VECTOR(11 DOWNTO 0);
	TYPE victory_image_type IS ARRAY (0 TO 39, 0 TO 311) OF STD_LOGIC_VECTOR(11 DOWNTO 0);
	
	-- Constant definition for the snake image
	CONSTANT snake_image : image_type := (
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"2B4", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000")
	);
	
	-- Constant definition for the food image
	CONSTANT food_image : image_type := (
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"000", X"000", X"000", X"000", X"000", X"000", X"FC0", X"000", X"000", X"000", X"000", X"000", X"000", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000", X"FC0", X"FC0", X"000", X"000", X"000", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"000", X"000", X"000", X"000", X"000", X"000", X"FC0", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000", X"000", X"000", X"000", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"FC0", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000")
	);
	
	-- Constant definition for the victory image
	CONSTANT victory_image : victory_image_type := (
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12")
	);
	
	-- Constant definition for the game over image
	CONSTANT gameOver_image : gameOver_image_type := (
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12")
	);
	
	-- Constant definition for the lives image
	CONSTANT live_image : image_type := (
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"E12", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"E12", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000"),
		(X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000", X"000")
	);

END PACKAGE snake_pkg;

PACKAGE BODY snake_pkg IS
END PACKAGE BODY snake_pkg;
